// Include file for sv_include_semicolon1 test
`define INCLUDED_VALUE 100
